//---------------------------------------------------------------------------
// Wishbone General Pupose IO Component
//
//     0x00	
//     
//     0x14     number   (read/write)
//    
//
//---------------------------------------------------------------------------

module wb_BCD (
	input              clk,
	input              reset,
	// Wishbone interface
	input              wb_stb_i,
	input              wb_cyc_i,
	output             wb_ack_o,
	input              wb_we_i,
	input       [31:0] wb_adr_i,
	input        [3:0] wb_sel_i,
	input       [31:0] wb_dat_i,
	output reg  [31:0] wb_dat_o,
	output [6:0] seg_out,
	output [3:0] an_out
);

//---------------------------------------------------------------------------
// 
//---------------------------------------------------------------------------

wire [31:0] BCDcr = 32'b0;

wire [6:0] seg0;
wire [3:0] an0;
reg [3:0] dato1;
reg [3:0] dato2;
reg [3:0] dato3;
reg [3:0] dato4;

BCD bcd0 (
	.clk(clk),
	.dato1(dato1),
	.dato2(dato2),
	.dato3(dato3),
	.dato4(dato4),
	.seg(seg0),
	.an(an0)
);


// Wishbone
reg  ack;
assign wb_ack_o = wb_stb_i & wb_cyc_i & ack;

wire wb_rd = wb_stb_i & wb_cyc_i & ~wb_we_i;
wire wb_wr = wb_stb_i & wb_cyc_i &  wb_we_i;



always @(posedge clk)
begin
	if (reset) begin
		ack      <= 0;
dato1<=15;
dato2<=15;
dato3<=15;
dato4<=15;

		
	end else begin
		// Handle WISHBONE access
		ack    <= 0;

		if (wb_wr & ~ack ) begin // write cycle
			ack <= 1;

			case (wb_adr_i[3:2])
			2'b00: dato1 <= wb_dat_i[3:0];	//wb_dat_i		
			2'b01: dato2 <= wb_dat_i[3:0];			
			2'b10: dato3 <= wb_dat_i[3:0];			
			2'b11: dato4 <= wb_dat_i[3:0];			
			endcase
		end
	end
end


assign an_out = an0;
assign seg_out = seg0;


endmodule
